///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: MUX4
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: A, B, C, D (32-bit), S (2-bit)
reg[31:0] A;
reg[31:0] B;
reg[31:0] C;
reg[31:0] D;
reg[1:0] S;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: Y (32-bit)
wire[31:0] Y;
///////////////////////////////////////////////////////////////////////////////////

MUX4_32 myMUX(.A(A), .B(B), .C(C), .D(D), .S(S), .Y(Y));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: S=00
$display("Testing: S=00");
A=32767; B=16383; C=65535; D=2481; S=2'b00;  #10; 
verifyEqual32(Y, A);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=01
$display("Testing: S=01");
S=2'b01;  #10; 
verifyEqual32(Y, B);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=10
$display("Testing: S=10");
S=2'b10;  #10; 
verifyEqual32(Y, C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=11
$display("Testing: S=11");
S=2'b11;  #10; 
verifyEqual32(Y, D);
////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule